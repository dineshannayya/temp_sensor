module tempsenseInst_error (CLK_REF,
    DONE,
    RESET_COUNTERn,
    en,
    lc_out,
    out,
    outb,
    DOUT,
    SEL_CONV_TIME);
 input CLK_REF;
 output DONE;
 input RESET_COUNTERn;
 input en;
 output lc_out;
 output out;
 output outb;
 output [23:0] DOUT;
 input [3:0] SEL_CONV_TIME;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire \temp_analog_0.n1 ;
 wire \temp_analog_0.n2 ;
 wire \temp_analog_0.n3 ;
 wire \temp_analog_0.n4 ;
 wire \temp_analog_0.n5 ;
 wire \temp_analog_0.n6 ;
 wire \temp_analog_0.n7 ;
 wire \temp_analog_0.nx2 ;
 wire \temp_analog_1.VIN ;
 wire \temp_analog_1.async_counter_0.WAKE ;
 wire \temp_analog_1.async_counter_0.WAKE_pre ;
 wire \temp_analog_1.async_counter_0.clk_ref_in ;
 wire \temp_analog_1.async_counter_0.clk_sens_in ;
 wire \temp_analog_1.async_counter_0.div_r[0] ;
 wire \temp_analog_1.async_counter_0.div_r[10] ;
 wire \temp_analog_1.async_counter_0.div_r[11] ;
 wire \temp_analog_1.async_counter_0.div_r[12] ;
 wire \temp_analog_1.async_counter_0.div_r[13] ;
 wire \temp_analog_1.async_counter_0.div_r[14] ;
 wire \temp_analog_1.async_counter_0.div_r[15] ;
 wire \temp_analog_1.async_counter_0.div_r[16] ;
 wire \temp_analog_1.async_counter_0.div_r[17] ;
 wire \temp_analog_1.async_counter_0.div_r[18] ;
 wire \temp_analog_1.async_counter_0.div_r[19] ;
 wire \temp_analog_1.async_counter_0.div_r[1] ;
 wire \temp_analog_1.async_counter_0.div_r[20] ;
 wire \temp_analog_1.async_counter_0.div_r[2] ;
 wire \temp_analog_1.async_counter_0.div_r[3] ;
 wire \temp_analog_1.async_counter_0.div_r[4] ;
 wire \temp_analog_1.async_counter_0.div_r[5] ;
 wire \temp_analog_1.async_counter_0.div_r[6] ;
 wire \temp_analog_1.async_counter_0.div_r[7] ;
 wire \temp_analog_1.async_counter_0.div_r[8] ;
 wire \temp_analog_1.async_counter_0.div_r[9] ;
 wire \temp_analog_1.async_counter_0.div_s[0] ;
 wire \temp_analog_1.async_counter_0.div_s[10] ;
 wire \temp_analog_1.async_counter_0.div_s[11] ;
 wire \temp_analog_1.async_counter_0.div_s[12] ;
 wire \temp_analog_1.async_counter_0.div_s[13] ;
 wire \temp_analog_1.async_counter_0.div_s[14] ;
 wire \temp_analog_1.async_counter_0.div_s[15] ;
 wire \temp_analog_1.async_counter_0.div_s[16] ;
 wire \temp_analog_1.async_counter_0.div_s[17] ;
 wire \temp_analog_1.async_counter_0.div_s[18] ;
 wire \temp_analog_1.async_counter_0.div_s[19] ;
 wire \temp_analog_1.async_counter_0.div_s[1] ;
 wire \temp_analog_1.async_counter_0.div_s[20] ;
 wire \temp_analog_1.async_counter_0.div_s[21] ;
 wire \temp_analog_1.async_counter_0.div_s[22] ;
 wire \temp_analog_1.async_counter_0.div_s[23] ;
 wire \temp_analog_1.async_counter_0.div_s[2] ;
 wire \temp_analog_1.async_counter_0.div_s[3] ;
 wire \temp_analog_1.async_counter_0.div_s[4] ;
 wire \temp_analog_1.async_counter_0.div_s[5] ;
 wire \temp_analog_1.async_counter_0.div_s[6] ;
 wire \temp_analog_1.async_counter_0.div_s[7] ;
 wire \temp_analog_1.async_counter_0.div_s[8] ;
 wire \temp_analog_1.async_counter_0.div_s[9] ;

 sky130_fd_sc_hd__fill_2 FILLER_0_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_0_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_0_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_0_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_0_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_0_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_0_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_10_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_10_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_10_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_10_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_10_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_10_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_10_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_10_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_10_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_10_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_10_86 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_11_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_11_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_11_171 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_11_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_11_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_11_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_230 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_11_242 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_11_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_11_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_11_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_11_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_11_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_12_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_12_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_12_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_12_170 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_182 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_12_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_12_198 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_12_202 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_12_211 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_12_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_12_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_12_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_12_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_12_86 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_13_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_13_143 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_13_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_13_172 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_13_183 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_13_191 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_13_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_216 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_228 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_13_240 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_13_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_13_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_13_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_13_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_13_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_13_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_14_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_14_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_14_155 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_14_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_14_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_173 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_14_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_14_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_14_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_14_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_14_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_14_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_14_89 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_14_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_15_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_15_143 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_171 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_15_183 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_15_191 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_15_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_15_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_15_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_15_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_15_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_15_76 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_15_80 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_15_87 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_15_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_15_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_16_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_16_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_16_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_16_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_16_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_16_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_16_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_16_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_16_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_16_73 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_16_80 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_16_87 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_16_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_16_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_17_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_17_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_17_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_17_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_17_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_17_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_17_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_18_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_18_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_18_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_18_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_18_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_18_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_18_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_18_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_19_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_19_170 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_19_182 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_19_190 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_19_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_19_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_19_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_19_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_19_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_19_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_19_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_1_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_1_186 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_1_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_1_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_1_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_1_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_20_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_20_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_20_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_20_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_20_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_20_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_175 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_21_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_21_191 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_21_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_21_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_21_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_21_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_22_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_22_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_22_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_22_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_22_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_22_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_23_108 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_23_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_133 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_138 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_23_164 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_23_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_23_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_23_208 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_23_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_23_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_23_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_23_37 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_23_45 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_54 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_23_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_23_61 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_23_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_23_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_23_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_23_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_108 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_120 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_24_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_24_188 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_232 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_24_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_24_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_24_58 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_24_68 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_24_75 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_82 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_24_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_25_107 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_25_111 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_137 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_149 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_25_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_25_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_25_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_25_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_25_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_25_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_25_61 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_25_95 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_109 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_121 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_26_133 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_26_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_239 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_26_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_26_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_26_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_26_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_27_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_27_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_27_121 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_128 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_140 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_152 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_27_164 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_27_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_27_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_27_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_27_93 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_28_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_28_111 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_28_136 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_28_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_28_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_28_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_28_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_28_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_28_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_28_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_29_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_29_109 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_29_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_120 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_132 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_29_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_29_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_29_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_29_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_29_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_29_93 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_2_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_2_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_2_154 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_2_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_2_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_2_173 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_2_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_2_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_2_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_2_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_2_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_2_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_2_243 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_2_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_117 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_30_129 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_30_137 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_30_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_30_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_30_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_30_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_30_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_30_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_30_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_30_93 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_31_102 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_31_110 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_137 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_149 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_31_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_31_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_31_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_31_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_31_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_31_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_31_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_31_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_31_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_109 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_121 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_32_133 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_153 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_32_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_32_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_32_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_32_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_32_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_32_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_32_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_32_66 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_32_73 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_32_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_32_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_33_108 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_33_137 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_33_145 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_33_150 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_33_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_33_166 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_33_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_33_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_33_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_33_223 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_33_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_33_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_33_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_33_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_33_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_109 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_121 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_34_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_176 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_192 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_34_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_34_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_34_45 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_49 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_34_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_34_92 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_34_99 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_35_109 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_35_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_35_118 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_35_124 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_128 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_135 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_142 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_35_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_152 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_163 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_35_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_192 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_35_199 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_35_206 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_35_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_35_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_35_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_35_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_35_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_35_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_35_54 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_35_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_35_80 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_36_119 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_36_127 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_131 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_36_138 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_36_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_168 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_36_172 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_36_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_36_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_212 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_224 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_236 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_248 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_36_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_36_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_36_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_36_82 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_36_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_36_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_37_101 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_37_110 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_37_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_37_136 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_37_140 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_37_162 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_37_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_37_178 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_37_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_37_215 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_37_222 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_37_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_37_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_37_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_37_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_37_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_37_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_37_76 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_38_106 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_38_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_138 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_38_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_38_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_38_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_239 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_38_251 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_38_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_38_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_38_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_61 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_38_66 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_38_73 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_38_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_38_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_38_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_38_99 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_103 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_39_110 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_39_117 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_125 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_39_150 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_39_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_39_166 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_39_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_39_181 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_39_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_209 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_39_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_230 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_242 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_39_254 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_39_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_39_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_39_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_89 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_39_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_3_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_3_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_3_172 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_3_184 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_3_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_3_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_3_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_3_212 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_3_216 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_3_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_3_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_3_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_3_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_3_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_103 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_40_138 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_40_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_187 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_40_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_40_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_40_227 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_234 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_40_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_40_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_40_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_40_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_40_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_40_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_40_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_110 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_113 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_136 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_41_141 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_154 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_166 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_169 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_174 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_185 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_194 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_197 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_206 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_41_220 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_225 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_237 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_41_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_41_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_41_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_41_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_41_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_41_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_41_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_4_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_4_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_4_154 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_4_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_4_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_4_188 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_4_196 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_4_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_4_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_4_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_4_252 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_5_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_5_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_5_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_5_158 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_5_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_5_173 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_5_180 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_5_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_5_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_5_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_5_244 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_5_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_6_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_6_154 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_6_161 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_6_188 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_6_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_206 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_218 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_226 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_6_238 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_6_246 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_6_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_6_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_6_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 FILLER_6_86 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_6_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_7_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_7_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_7_151 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_176 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_7_188 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_7_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_7_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_7_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_7_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_7_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_7_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_7_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_8_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_144 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_8_156 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_165 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_177 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_189 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_201 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_8_213 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_8_219 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_221 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_233 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_8_245 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_8_253 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_8_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_8_86 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_2 FILLER_9_139 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_147 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_159 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_171 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_9_183 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_9_191 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_193 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_205 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_217 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_229 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_9_241 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_9_247 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_6 FILLER_9_249 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_ef_sc_hd__decap_12 FILLER_9_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_4 FILLER_9_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__fill_1 FILLER_9_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_8 FILLER_9_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(VSS),
    .VPWR(VIN));
 sky130_fd_sc_hd__inv_2 _108_ (.A(\temp_analog_1.async_counter_0.div_r[5] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _109_ (.A(SEL_CONV_TIME[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _110_ (.A(\temp_analog_1.async_counter_0.div_r[20] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(\temp_analog_1.async_counter_0.div_r[19] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _112_ (.A(\temp_analog_1.async_counter_0.div_r[18] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _113_ (.A(\temp_analog_1.async_counter_0.div_r[17] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _114_ (.A(\temp_analog_1.async_counter_0.div_r[16] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _115_ (.A(\temp_analog_1.async_counter_0.div_r[15] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _116_ (.A(\temp_analog_1.async_counter_0.div_r[14] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(\temp_analog_1.async_counter_0.div_r[13] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _118_ (.A(\temp_analog_1.async_counter_0.div_r[12] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _119_ (.A(\temp_analog_1.async_counter_0.div_r[11] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _120_ (.A(\temp_analog_1.async_counter_0.div_r[10] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _121_ (.A(\temp_analog_1.async_counter_0.div_r[9] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _122_ (.A(\temp_analog_1.async_counter_0.div_r[8] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _123_ (.A(\temp_analog_1.async_counter_0.div_r[7] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _124_ (.A(\temp_analog_1.async_counter_0.div_r[6] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _125_ (.A(\temp_analog_1.async_counter_0.div_s[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _126_ (.A(\temp_analog_1.async_counter_0.div_s[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _127_ (.A(\temp_analog_1.async_counter_0.div_s[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _128_ (.A(\temp_analog_1.async_counter_0.div_s[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _129_ (.A(\temp_analog_1.async_counter_0.div_s[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _130_ (.A(\temp_analog_1.async_counter_0.div_s[5] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _131_ (.A(\temp_analog_1.async_counter_0.div_s[6] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _132_ (.A(\temp_analog_1.async_counter_0.div_s[7] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _133_ (.A(\temp_analog_1.async_counter_0.div_s[8] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _134_ (.A(\temp_analog_1.async_counter_0.div_s[9] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(\temp_analog_1.async_counter_0.div_s[10] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _136_ (.A(\temp_analog_1.async_counter_0.div_s[11] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _137_ (.A(\temp_analog_1.async_counter_0.div_s[12] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _138_ (.A(\temp_analog_1.async_counter_0.div_s[13] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _139_ (.A(\temp_analog_1.async_counter_0.div_s[14] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _140_ (.A(\temp_analog_1.async_counter_0.div_s[15] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _141_ (.A(\temp_analog_1.async_counter_0.div_s[16] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _142_ (.A(\temp_analog_1.async_counter_0.div_s[17] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _143_ (.A(\temp_analog_1.async_counter_0.div_s[18] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _144_ (.A(\temp_analog_1.async_counter_0.div_s[19] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _145_ (.A(\temp_analog_1.async_counter_0.div_s[20] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _146_ (.A(\temp_analog_1.async_counter_0.div_s[21] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _147_ (.A(\temp_analog_1.async_counter_0.div_s[22] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _148_ (.A(\temp_analog_1.async_counter_0.div_s[23] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _149_ (.A(\temp_analog_1.async_counter_0.div_r[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _150_ (.A(\temp_analog_1.async_counter_0.div_r[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _151_ (.A(\temp_analog_1.async_counter_0.div_r[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _152_ (.A(\temp_analog_1.async_counter_0.div_r[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _153_ (.A(\temp_analog_1.async_counter_0.div_r[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_004_));
 sky130_fd_sc_hd__or3b_2 _154_ (.A(SEL_CONV_TIME[0]),
    .B(\temp_analog_1.async_counter_0.div_r[11] ),
    .C_N(SEL_CONV_TIME[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_089_));
 sky130_fd_sc_hd__nand2b_2 _155_ (.A_N(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_2 _156_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_091_));
 sky130_fd_sc_hd__or3_2 _157_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(\temp_analog_1.async_counter_0.div_r[9] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_092_));
 sky130_fd_sc_hd__o221a_2 _158_ (.A1(\temp_analog_1.async_counter_0.div_r[10] ),
    .A2(_090_),
    .B1(_091_),
    .B2(\temp_analog_1.async_counter_0.div_r[12] ),
    .C1(_092_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_093_));
 sky130_fd_sc_hd__and3b_2 _159_ (.A_N(SEL_CONV_TIME[3]),
    .B(_089_),
    .C(_093_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_094_));
 sky130_fd_sc_hd__or3b_2 _160_ (.A(SEL_CONV_TIME[0]),
    .B(\temp_analog_1.async_counter_0.div_r[19] ),
    .C_N(SEL_CONV_TIME[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_095_));
 sky130_fd_sc_hd__or3_2 _161_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(\temp_analog_1.async_counter_0.div_r[17] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_096_));
 sky130_fd_sc_hd__o221a_2 _162_ (.A1(\temp_analog_1.async_counter_0.div_r[18] ),
    .A2(_090_),
    .B1(_091_),
    .B2(\temp_analog_1.async_counter_0.div_r[20] ),
    .C1(_096_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_097_));
 sky130_fd_sc_hd__a31o_2 _163_ (.A1(SEL_CONV_TIME[3]),
    .A2(_095_),
    .A3(_097_),
    .B1(_088_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_098_));
 sky130_fd_sc_hd__mux4_2 _164_ (.A0(\temp_analog_1.async_counter_0.div_r[5] ),
    .A1(\temp_analog_1.async_counter_0.div_r[7] ),
    .A2(\temp_analog_1.async_counter_0.div_r[6] ),
    .A3(\temp_analog_1.async_counter_0.div_r[8] ),
    .S0(SEL_CONV_TIME[1]),
    .S1(SEL_CONV_TIME[0]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_099_));
 sky130_fd_sc_hd__nand2b_2 _165_ (.A_N(SEL_CONV_TIME[3]),
    .B(_099_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_100_));
 sky130_fd_sc_hd__or2_2 _166_ (.A(\temp_analog_1.async_counter_0.div_r[14] ),
    .B(_090_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_101_));
 sky130_fd_sc_hd__or3b_2 _167_ (.A(SEL_CONV_TIME[0]),
    .B(\temp_analog_1.async_counter_0.div_r[15] ),
    .C_N(SEL_CONV_TIME[1]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_102_));
 sky130_fd_sc_hd__or3_2 _168_ (.A(SEL_CONV_TIME[1]),
    .B(SEL_CONV_TIME[0]),
    .C(\temp_analog_1.async_counter_0.div_r[13] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_103_));
 sky130_fd_sc_hd__o2111a_2 _169_ (.A1(\temp_analog_1.async_counter_0.div_r[16] ),
    .A2(_091_),
    .B1(_102_),
    .C1(_103_),
    .D1(SEL_CONV_TIME[3]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_104_));
 sky130_fd_sc_hd__a21oi_2 _170_ (.A1(_101_),
    .A2(_104_),
    .B1(SEL_CONV_TIME[2]),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_105_));
 sky130_fd_sc_hd__o2bb2a_2 _171_ (.A1_N(_105_),
    .A2_N(_100_),
    .B1(_098_),
    .B2(_094_),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DONE));
 sky130_fd_sc_hd__and3b_2 _172_ (.A_N(DONE),
    .B(CLK_REF),
    .C(\temp_analog_1.async_counter_0.WAKE ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(\temp_analog_1.async_counter_0.clk_ref_in ));
 sky130_fd_sc_hd__and3b_2 _173_ (.A_N(DONE),
    .B(lc_out),
    .C(\temp_analog_1.async_counter_0.WAKE_pre ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(\temp_analog_1.async_counter_0.clk_sens_in ));
 sky130_fd_sc_hd__and2_2 _174_ (.A(\temp_analog_1.async_counter_0.div_s[0] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[0]));
 sky130_fd_sc_hd__and2_2 _175_ (.A(\temp_analog_1.async_counter_0.div_s[1] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[1]));
 sky130_fd_sc_hd__and2_2 _176_ (.A(\temp_analog_1.async_counter_0.div_s[2] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[2]));
 sky130_fd_sc_hd__and2_2 _177_ (.A(\temp_analog_1.async_counter_0.div_s[3] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[3]));
 sky130_fd_sc_hd__and2_2 _178_ (.A(\temp_analog_1.async_counter_0.div_s[4] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[4]));
 sky130_fd_sc_hd__and2_2 _179_ (.A(\temp_analog_1.async_counter_0.div_s[5] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[5]));
 sky130_fd_sc_hd__and2_2 _180_ (.A(\temp_analog_1.async_counter_0.div_s[6] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[6]));
 sky130_fd_sc_hd__and2_2 _181_ (.A(\temp_analog_1.async_counter_0.div_s[7] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[7]));
 sky130_fd_sc_hd__and2_2 _182_ (.A(\temp_analog_1.async_counter_0.div_s[8] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[8]));
 sky130_fd_sc_hd__and2_2 _183_ (.A(\temp_analog_1.async_counter_0.div_s[9] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[9]));
 sky130_fd_sc_hd__and2_2 _184_ (.A(\temp_analog_1.async_counter_0.div_s[10] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[10]));
 sky130_fd_sc_hd__and2_2 _185_ (.A(\temp_analog_1.async_counter_0.div_s[11] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[11]));
 sky130_fd_sc_hd__and2_2 _186_ (.A(\temp_analog_1.async_counter_0.div_s[12] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[12]));
 sky130_fd_sc_hd__and2_2 _187_ (.A(\temp_analog_1.async_counter_0.div_s[13] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[13]));
 sky130_fd_sc_hd__and2_2 _188_ (.A(\temp_analog_1.async_counter_0.div_s[14] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[14]));
 sky130_fd_sc_hd__and2_2 _189_ (.A(\temp_analog_1.async_counter_0.div_s[15] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[15]));
 sky130_fd_sc_hd__and2_2 _190_ (.A(\temp_analog_1.async_counter_0.div_s[16] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[16]));
 sky130_fd_sc_hd__and2_2 _191_ (.A(\temp_analog_1.async_counter_0.div_s[17] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[17]));
 sky130_fd_sc_hd__and2_2 _192_ (.A(\temp_analog_1.async_counter_0.div_s[18] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[18]));
 sky130_fd_sc_hd__and2_2 _193_ (.A(\temp_analog_1.async_counter_0.div_s[19] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[19]));
 sky130_fd_sc_hd__and2_2 _194_ (.A(\temp_analog_1.async_counter_0.div_s[20] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[20]));
 sky130_fd_sc_hd__and2_2 _195_ (.A(\temp_analog_1.async_counter_0.div_s[21] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[21]));
 sky130_fd_sc_hd__and2_2 _196_ (.A(\temp_analog_1.async_counter_0.div_s[22] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[22]));
 sky130_fd_sc_hd__and2_2 _197_ (.A(\temp_analog_1.async_counter_0.div_s[23] ),
    .B(DONE),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(DOUT[23]));
 sky130_fd_sc_hd__or2_2 _198_ (.A(\temp_analog_1.async_counter_0.WAKE ),
    .B(\temp_analog_1.async_counter_0.WAKE_pre ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .X(_072_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(\temp_analog_1.async_counter_0.div_r[19] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(\temp_analog_1.async_counter_0.div_r[18] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(\temp_analog_1.async_counter_0.div_r[17] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _202_ (.A(\temp_analog_1.async_counter_0.div_r[16] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(\temp_analog_1.async_counter_0.div_r[15] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(\temp_analog_1.async_counter_0.div_r[14] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(\temp_analog_1.async_counter_0.div_r[13] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(\temp_analog_1.async_counter_0.div_r[12] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(\temp_analog_1.async_counter_0.div_r[11] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(\temp_analog_1.async_counter_0.div_r[10] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(\temp_analog_1.async_counter_0.div_r[9] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _210_ (.A(\temp_analog_1.async_counter_0.div_r[8] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _211_ (.A(\temp_analog_1.async_counter_0.div_r[7] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _212_ (.A(\temp_analog_1.async_counter_0.div_r[6] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _213_ (.A(\temp_analog_1.async_counter_0.div_r[5] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(\temp_analog_1.async_counter_0.div_r[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _215_ (.A(\temp_analog_1.async_counter_0.div_r[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _216_ (.A(\temp_analog_1.async_counter_0.div_r[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _217_ (.A(\temp_analog_1.async_counter_0.div_r[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(\temp_analog_1.async_counter_0.div_r[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _219_ (.A(\temp_analog_1.async_counter_0.div_s[22] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(\temp_analog_1.async_counter_0.div_s[21] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _221_ (.A(\temp_analog_1.async_counter_0.div_s[20] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(\temp_analog_1.async_counter_0.div_s[19] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _223_ (.A(\temp_analog_1.async_counter_0.div_s[18] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _224_ (.A(\temp_analog_1.async_counter_0.div_s[17] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _225_ (.A(\temp_analog_1.async_counter_0.div_s[16] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_065_));
 sky130_fd_sc_hd__inv_2 _226_ (.A(\temp_analog_1.async_counter_0.div_s[15] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _227_ (.A(\temp_analog_1.async_counter_0.div_s[14] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(\temp_analog_1.async_counter_0.div_s[13] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _229_ (.A(\temp_analog_1.async_counter_0.div_s[12] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _230_ (.A(\temp_analog_1.async_counter_0.div_s[11] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _231_ (.A(\temp_analog_1.async_counter_0.div_s[10] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _232_ (.A(\temp_analog_1.async_counter_0.div_s[9] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(\temp_analog_1.async_counter_0.div_s[8] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _234_ (.A(\temp_analog_1.async_counter_0.div_s[7] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _235_ (.A(\temp_analog_1.async_counter_0.div_s[6] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _236_ (.A(\temp_analog_1.async_counter_0.div_s[5] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(\temp_analog_1.async_counter_0.div_s[4] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(\temp_analog_1.async_counter_0.div_s[3] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\temp_analog_1.async_counter_0.div_s[2] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(\temp_analog_1.async_counter_0.div_s[1] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(\temp_analog_1.async_counter_0.div_s[0] ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(_038_));
 sky130_fd_sc_hd__dfrtp_2 _242_ (.CLK(CLK_REF),
    .D(_072_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.WAKE ));
 sky130_fd_sc_hd__dfrtp_2 _243_ (.CLK(CLK_REF),
    .D(_106_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.WAKE_pre ));
 sky130_fd_sc_hd__dfrtp_2 _244_ (.CLK(_039_),
    .D(_073_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[20] ));
 sky130_fd_sc_hd__dfrtp_2 _245_ (.CLK(_040_),
    .D(_079_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[19] ));
 sky130_fd_sc_hd__dfrtp_2 _246_ (.CLK(_041_),
    .D(_080_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[18] ));
 sky130_fd_sc_hd__dfrtp_2 _247_ (.CLK(_042_),
    .D(_081_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[17] ));
 sky130_fd_sc_hd__dfrtp_2 _248_ (.CLK(_043_),
    .D(_082_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[16] ));
 sky130_fd_sc_hd__dfrtp_2 _249_ (.CLK(_044_),
    .D(_083_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[15] ));
 sky130_fd_sc_hd__dfrtp_2 _250_ (.CLK(_045_),
    .D(_084_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[14] ));
 sky130_fd_sc_hd__dfrtp_2 _251_ (.CLK(_046_),
    .D(_085_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[13] ));
 sky130_fd_sc_hd__dfrtp_2 _252_ (.CLK(_047_),
    .D(_086_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[12] ));
 sky130_fd_sc_hd__dfrtp_2 _253_ (.CLK(_048_),
    .D(_087_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[11] ));
 sky130_fd_sc_hd__dfrtp_2 _254_ (.CLK(_049_),
    .D(_074_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[10] ));
 sky130_fd_sc_hd__dfrtp_2 _255_ (.CLK(_050_),
    .D(_075_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[9] ));
 sky130_fd_sc_hd__dfrtp_2 _256_ (.CLK(_051_),
    .D(_076_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[8] ));
 sky130_fd_sc_hd__dfrtp_2 _257_ (.CLK(_052_),
    .D(_077_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[7] ));
 sky130_fd_sc_hd__dfrtp_2 _258_ (.CLK(_053_),
    .D(_078_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[6] ));
 sky130_fd_sc_hd__dfrtp_2 _259_ (.CLK(_054_),
    .D(_107_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[5] ));
 sky130_fd_sc_hd__dfrtp_2 _260_ (.CLK(_055_),
    .D(_004_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[4] ));
 sky130_fd_sc_hd__dfrtp_2 _261_ (.CLK(_056_),
    .D(_003_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[3] ));
 sky130_fd_sc_hd__dfrtp_2 _262_ (.CLK(_057_),
    .D(_002_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[2] ));
 sky130_fd_sc_hd__dfrtp_2 _263_ (.CLK(_058_),
    .D(_001_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[1] ));
 sky130_fd_sc_hd__dfrtp_2 _264_ (.CLK(_059_),
    .D(_020_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[23] ));
 sky130_fd_sc_hd__dfrtp_2 _265_ (.CLK(_060_),
    .D(_019_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[22] ));
 sky130_fd_sc_hd__dfrtp_2 _266_ (.CLK(_061_),
    .D(_018_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[21] ));
 sky130_fd_sc_hd__dfrtp_2 _267_ (.CLK(_062_),
    .D(_017_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[20] ));
 sky130_fd_sc_hd__dfrtp_2 _268_ (.CLK(_063_),
    .D(_015_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[19] ));
 sky130_fd_sc_hd__dfrtp_2 _269_ (.CLK(_064_),
    .D(_014_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[18] ));
 sky130_fd_sc_hd__dfrtp_2 _270_ (.CLK(_065_),
    .D(_013_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[17] ));
 sky130_fd_sc_hd__dfrtp_2 _271_ (.CLK(_066_),
    .D(_012_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[16] ));
 sky130_fd_sc_hd__dfrtp_2 _272_ (.CLK(_067_),
    .D(_011_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[15] ));
 sky130_fd_sc_hd__dfrtp_2 _273_ (.CLK(_068_),
    .D(_010_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[14] ));
 sky130_fd_sc_hd__dfrtp_2 _274_ (.CLK(_069_),
    .D(_009_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[13] ));
 sky130_fd_sc_hd__dfrtp_2 _275_ (.CLK(_070_),
    .D(_008_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[12] ));
 sky130_fd_sc_hd__dfrtp_2 _276_ (.CLK(_071_),
    .D(_007_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[11] ));
 sky130_fd_sc_hd__dfrtp_2 _277_ (.CLK(_029_),
    .D(_006_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[10] ));
 sky130_fd_sc_hd__dfrtp_2 _278_ (.CLK(_030_),
    .D(_028_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[9] ));
 sky130_fd_sc_hd__dfrtp_2 _279_ (.CLK(_031_),
    .D(_027_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[8] ));
 sky130_fd_sc_hd__dfrtp_2 _280_ (.CLK(_032_),
    .D(_026_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[7] ));
 sky130_fd_sc_hd__dfrtp_2 _281_ (.CLK(_033_),
    .D(_025_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[6] ));
 sky130_fd_sc_hd__dfrtp_2 _282_ (.CLK(_034_),
    .D(_024_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[5] ));
 sky130_fd_sc_hd__dfrtp_2 _283_ (.CLK(_035_),
    .D(_023_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[4] ));
 sky130_fd_sc_hd__dfrtp_2 _284_ (.CLK(_036_),
    .D(_022_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[3] ));
 sky130_fd_sc_hd__dfrtp_2 _285_ (.CLK(_037_),
    .D(_021_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[2] ));
 sky130_fd_sc_hd__dfrtp_2 _286_ (.CLK(_038_),
    .D(_016_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[1] ));
 sky130_fd_sc_hd__dfrtp_2 _287_ (.CLK(\temp_analog_1.async_counter_0.clk_ref_in ),
    .D(_000_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_r[0] ));
 sky130_fd_sc_hd__dfrtp_2 _288_ (.CLK(\temp_analog_1.async_counter_0.clk_sens_in ),
    .D(_005_),
    .RESET_B(RESET_COUNTERn),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Q(\temp_analog_1.async_counter_0.div_s[0] ));
 sky130_fd_sc_hd__conb_1 _289_ (.VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .HI(_106_));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_0  (.A(\temp_analog_0.n1 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n2 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_1  (.A(\temp_analog_0.n2 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n3 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_2  (.A(\temp_analog_0.n3 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n4 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_3  (.A(\temp_analog_0.n4 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n5 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_4  (.A(\temp_analog_0.n5 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n6 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_5  (.A(\temp_analog_0.n6 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n7 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m1  (.A(\temp_analog_0.n7 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(out));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m2  (.A(\temp_analog_0.n7 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.nx2 ));
 sky130_fd_sc_hd__inv_1 \temp_analog_0.a_inv_m3  (.A(\temp_analog_0.nx2 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(outb));
 sky130_fd_sc_hd__nand2_1 \temp_analog_0.a_nand_0  (.A(en),
    .B(\temp_analog_0.n7 ),
    .VGND(VSS),
    .VNB(VSS),
    .VPB(VIN),
    .VPWR(VIN),
    .Y(\temp_analog_0.n1 ));
 HEADER \temp_analog_1.a_header_0  (.VIN(\temp_analog_1.VIN ),
    .VNB(VSS),
    .VGND(VSS),
    .VPWR(VIN));
 HEADER \temp_analog_1.a_header_1  (.VIN(\temp_analog_1.VIN ),
    .VNB(VSS),
    .VGND(VSS),
    .VPWR(VIN));
 HEADER \temp_analog_1.a_header_2  (.VIN(\temp_analog_1.VIN ),
    .VNB(VSS),
    .VGND(VSS),
    .VPWR(VIN));
 SLC \temp_analog_1.a_lc_0  (.IN(out),
    .INB(outb),
    .VGND(VSS),
    .VNB(VSS),
    .VOUT(lc_out),
    .VPB(VIN),
    .VPWR(VIN));
endmodule
